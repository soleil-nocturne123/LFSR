/*
	AUTHOR: PHAN HOAI HUONG NGUYEN
	DESCRIPTION: APPLICATION LOGIC MODULE OF THE AFU
*/